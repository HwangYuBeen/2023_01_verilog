library verilog;
use verilog.vl_types.all;
entity AND_gate is
    port(
        din             : in     vl_logic;
        dout            : out    vl_logic
    );
end AND_gate;
